`ifndef FAST_TRANSFER
`define FAST_TRANSFER

// transfer������: ��������, ��������, ������ 
typedef enum {DARK_CONTIG, BRIGHT_CONTIG, NON_CONTIG} fast_trans_kind;

// DARK_CONTIG
class dc_trans;
    

endclass




`endif 